

module Pack (
  // Управляющие сигналы
  input i_clk,
  input i_reset,
  // Входные данные
  input i_data,
  input i_valid,
  // Выходные данные
  output o_data,
  output reg o_valid
);

endmodule